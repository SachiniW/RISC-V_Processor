`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/03/2021 10:29:06 AM
// Design Name: 
// Module Name: InstMemory.v
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module InstMemory (
    input [31:0] PC,
    output [31:0] INST  
);
    
reg [31:0]  I_MEM   [0:256];

initial begin

    I_MEM[0] = 32'h02b1c393;    //xori x3 -> x7    0000  0010  1011,  0001  1,100, 0011  1,001 0011
    I_MEM[1] = 32'h00c3e793;    //ori  x7 -> x15   0000  0000  1100,  0011  1,110, 0111  1,001 0011
    I_MEM[2] = 32'h0317f493;    //andi x15-> x9    0000  0011  0001,  0111  1,111, 0100  1,001 0011
    I_MEM[3] = 32'h00748233;    //add  x9,x7->x4   0000  000,0 0111,  0100  1,000, 0010  0,011 0011
    I_MEM[4] = 32'h409208b3;    //sub  x4,x9->x17  0100  000,0 1001,  0010  0,000, 1000  1,011 0011
    I_MEM[5] = 32'h004792b3;    //sll  x15,x4->x5  0000  000,0 0100,  0111  1,001, 0010  1,011 0011
    I_MEM[6] = 32'h0034a783;    //lw mem[36]-> x15 0000  0000  0011,  0100  1,010, 0111  1,000 0011
    I_MEM[7] = 32'h01000f6f;    //jal->[44],rd=x30 0,000 0001  000,0, 0000  0,000, 1111  0,110 1111 //jump [28+16]
    I_MEM[8] = 32'h0034a203;    //lw mem[36]-> x4  0000  0000  0011,  0100  1,010, 0010  0,000 0011 <-bge target
    I_MEM[9] = 32'h0034a283;    //lw mem[36]-> x5  0000  0000  0011,  0100  1,010, 0010  1,000 0011
    I_MEM[10] = 32'h00924863;   //blt x4<x9->[56]  0000  000,0 1001,  0010  0,100, 1000  0,110 0011 //branch l [40+16]
    I_MEM[11] = 32'h00c3e793;   //ori  x7 -> x15   0000  0000  1100,  0011  1,110, 0111  1,001 0011 <- jal target
    I_MEM[12] = 32'hfffffa37;   //lui  rd -> x20   1111  1111  1111,  1111  1,111, 1010  0,011 0111 
    I_MEM[13] = 32'hff43d6e3;   //bge x7>x20->[32] 1111  111,1 0100,  0011  1,101, 0110  1,110 0011 //branch g [52-20]
    I_MEM[14] = 32'h0003e137;   //lui  rd -> x2    0000  0000  0000,  0011  1,110, 0001  0,011 0111  <- blt target
    

//    I_MEM[0] = 32'hfe010113;    //addi	sp,sp,-32
//    I_MEM[1] = 32'h02010413;   //addi	s0,sp,32
//    I_MEM[2] = 32'ha9478793;    //addi	a5,a5,-1388  # 0x10af8
//    I_MEM[3] = 32'h00178713;    //addi	a4,a5,1
//    I_MEM[4] = 32'h00f707b3;    //add	a5,a4,a5
//    I_MEM[5] = 32'h00271713;    //slli	a4,a4,0x2
//    I_MEM[6] = 32'h01045793;    //srli	a5,s0,0x10

end

assign INST = I_MEM[(PC>>2)];


endmodule



